-- ==============================================================
--  Lab 2 - VHDL Template
--  Descripci�n: Esqueleto de la entidad y arquitectura.
--  TODO: Completar descripci�n funcional del dise�o.
-- ==============================================================

-- TODO: A�adir librer�as necesarias.

entity uart_tx is
    port (
        -- TODO: A�adir puertos de entrada/salida.

    );
end entity uart_tx;

architecture RTL of uart_tx is

    -- ============================================================================
    -- DETECCI�N DE FLANCO DE SUBIDA DEL BOT�N
    -- ============================================================================
    -- TODO: Declarar constantes y tipos.
    -- TODO: Declarar se�ales internas.

    -- ============================================================================
    -- REGISTRO DE DESPLAZAMIENTO UART (Formato: 1 STOP + 8 DATOS + 1 START = 10 bits)
    -- ============================================================================
    -- TODO: Declarar constantes y tipos.
    -- TODO: Declarar se�ales internas.

    -- ============================================================================
    -- TEMPORIZADOR DE BIT (Controla duraci�n de cada bit a 19200 baud)
    -- Per�odo de bit = 100 MHz / 19200 = 5208 ciclos, limitado a 5207 = 13 bits
    -- ============================================================================
    -- TODO: Declarar constantes y tipos.
    -- TODO: Declarar se�ales internas.

begin

    -- ============================================================================
    -- DETECCI�N DE FLANCO DE SUBIDA DEL BOT�N
    -- ============================================================================
    -- ETAPA 1: SINCRONIZACI�N DEL BOT�N (2 registros de metaestabilidad)
    -- ETAPA 2: DEBOUNCING DEL BOT�N (Muestreo cada ~5 ms)
    -- ETAPA 3: DETECCI�N DE FLANCO DE SUBIDA

    -- TODO: Implementar el modelo separando parte combinacional de secuencial.


    -- ============================================================================
    -- REGISTRO DE DESPLAZAMIENTO UART
    -- ============================================================================

    -- TODO: Implementar el modelo separando parte combinacional de secuencial.

    -- ============================================================================
    -- TEMPORIZADOR DE BIT (timer para controlar duraci�n de cada bit)
    -- ============================================================================

    -- TODO: Implementar el modelo separando parte combinacional de secuencial.

    -- ============================================================================
    -- SALIDAS DEL M�DULO
    -- ============================================================================

    -- TODO: Asignar valores a los puertos de salida

end architecture;

